testbench.U_MUX
input_a
input_b
